Standard cell Simulation
* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

* instantiate the cell
Xcell A B VGND VNB VPB VPWR X sky130_fd_sc_hd__and2_0


